LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY mux3a1 IS
	PORT (
		A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		SEL_A : IN STD_LOGIC;
		SEL_B : IN STD_LOGIC;
		SEL_C : IN STD_LOGIC; 
		Y : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END mux3a1;

ARCHITECTURE Behavioral OF mux3a1 IS
BEGIN
	PROCESS (A, B, C, SEL_A, SEL_B, SEL_C)
	BEGIN
		IF SEL_A = '0' THEN
			Y <= A;
		ELSIF SEL_B = '0' THEN
			Y <= B;
		ELSIF SEL_C = '0' THEN
			Y <= C;
		ELSE
			-- Caso por defecto
			Y <= (OTHERS => 'X');
		END IF;
	END PROCESS;
END Behavioral;
